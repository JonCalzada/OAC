library ieee;
use ieee.std_logic_1164.all; 
use IEEE.std_logic_arith.all; 
use IEEE.std_logic_unsigned.all; 
entity memoria is 
port( dir: in std_logic_vector (3 downto 0); 
	data: out std_logic_vector (20 downto 0)); 
end memoria; 
architecture behavior of memoria is 
type mem is array (0 to 14) of std_logic_vector (20 downto 0);
signal s: mem;

begin 
	s(0)<="11"&"0"&"00"&"0000"&"000001"&"000001";
	s(1)<="00"&"1"&"01"&"0111"&"001111"&"001111";
	s(2)<="11"&"0"&"00"&"0000"&"000011"&"000011";
	s(3)<="11"&"0"&"00"&"0000"&"001010"&"001010";
	s(4)<="11"&"0"&"10"&"0000"&"010000"&"010000";
	s(5)<="01"&"1"&"01"&"1010"&"110010"&"010010";
	s(6)<="11"&"0"&"01"&"0010"&"001001"&"001001";
	s(7)<="10"&"1"&"11"&"0000"&"010001"&"010000";
	s(8)<="11"&"0"&"01"&"0001"&"100000"&"100000";
	s(9)<="10"&"0"&"11"&"0000"&"001010"&"101011";
	s(10)<="11"&"0"&"01"&"0000"&"001010"&"000000";
	s(11)<="11"&"0"&"10"&"0000"&"000100"&"000100";
	s(12)<="11"&"0"&"01"&"0000"&"000100"&"000100";
	s(13)<="11"&"0"&"01"&"0000"&"101000"&"101000";
	s(14)<="11"&"0"&"01"&"0000"&"010011"&"010011";
	
	process (dir)
		begin 
			data <= s(conv_integer(unsigned(dir)));
			end process;
		end behavior; 